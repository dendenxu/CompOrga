`timescale 1ns / 1ps

module multi_register_EN(
	EN,		// ʹ���źţ�����Ч��
	clk,		// ʱ���źţ������ش�����
	rst,		// ��λ�źţ�����Ч��
	data_in,	// ��������
	data_out	// �Ĵ������
);
	
	parameter N = 32;
	input  wire EN;
	input  wire clk, rst;
	input  wire [N - 1 : 0] data_in;
	output reg [N - 1 : 0] data_out;

	
	initial
		data_out = 0;

	always @(posedge clk or posedge rst)
		if (rst)
			data_out <= 0;
		else if (EN == 1'b1)
			data_out <= data_in;
		else
			data_out <= data_out;


endmodule
